conectix             �hevpc   Wi2k              ?   ���*�?I�9ހt�&��y�                                                                                                                                                                                                                                                                                                                                                                                                                                            cxsparse��������             �    ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                conectix             �hevpc   Wi2k              ?   ���*�?I�9ހt�&��y�                                                                                                                                                                                                                                                                                                                                                                                                                                            