conectix             ���vpc   Wi2k     �       �   �   ��티���އރZ�v_�                                                                                                                                                                                                                                                                                                                                                                                                                                            cxsparse��������                 ���s                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ����������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                conectix             ���vpc   Wi2k     �       �   �   ��티���އރZ�v_�                                                                                                                                                                                                                                                                                                                                                                                                                                            