conectix             �hXvpc   Wi2k              �   ��ﺅ?H�9ހt�&��y�                                                                                                                                                                                                                                                                                                                                                                                                                                            cxsparse��������             @    ���7                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                conectix             �hXvpc   Wi2k              �   ��ﺅ?H�9ހt�&��y�                                                                                                                                                                                                                                                                                                                                                                                                                                            